module dgldpc_shuffled_VNU
    (
        input  logic        [8 : 0] i_LOVNU                     ,
        input  logic                clk                         , 
        input  logic [0 : 3][5 : 0] i_data                      ,
        output logic [0 : 4][9 : 0] o_data      
    );    
    
endmodule